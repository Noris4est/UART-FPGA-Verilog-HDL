`timescale 1ns/1ps
module UART_TX_RX_MASSIV_MODULE_TB4
#(
	parameter UART_BAUD_RATE				=	9600,
   parameter CLOCK_FREQUENCY				=	38400,
   parameter PARITY							=	1,
   parameter NUM_OF_DATA_BITS_IN_PACK	=	8,
	parameter NUMBER_STOP_BITS				=	3,
	parameter TX_MASSIV_DEEP				=	2,
	parameter RX_MASSIV_DEEP				=	2,
	parameter RX_MASSIV_DEEP_LOG_2=$clog2(RX_MASSIV_DEEP),
	parameter TX_MASSIV_DEEP_LOG_2=$clog2(TX_MASSIV_DEEP)
);
localparam PERIOD_IN_CLOCK_NS=1000000000/CLOCK_FREQUENCY;
reg IN_CLOCK_1,	IN_CLOCK_2;
reg [NUM_OF_DATA_BITS_IN_PACK*TX_MASSIV_DEEP-1:0] IN_TX_DATA_MASSIV_1,	IN_TX_DATA_MASSIV_2;
reg [TX_MASSIV_DEEP_LOG_2:0] IN_TX_NUMBER_OF_PACKS_TO_SEND_1,	IN_TX_NUMBER_OF_PACKS_TO_SEND_2;
reg IN_TX_LAUNCH_1,IN_TX_LAUNCH_2;
reg IN_RX_CLEAR_BUFFER_1,IN_RX_CLEAR_BUFFER_2;

wire OUT_TX_ACTIVE_1,OUT_TX_ACTIVE_2;
wire OUT_TX_DONE_1,OUT_TX_DONE_2;
wire [NUM_OF_DATA_BITS_IN_PACK*RX_MASSIV_DEEP-1:0] OUT_RX_DATA_MASSIV_1,OUT_RX_DATA_MASSIV_2;
wire [RX_MASSIV_DEEP_LOG_2:0] OUT_RX_ERROR_1,OUT_RX_ERROR_2;
wire [RX_MASSIV_DEEP_LOG_2:0] OUT_RX_NUM_OF_DATA_PACKS_READY_1,OUT_RX_NUM_OF_DATA_PACKS_READY_2;


UART_TX_RX_MASSIV_MODULE
#(
	.UART_BAUD_RATE(UART_BAUD_RATE),
	.CLOCK_FREQUENCY(CLOCK_FREQUENCY),
	.PARITY(PARITY),
	.NUM_OF_DATA_BITS_IN_PACK(NUM_OF_DATA_BITS_IN_PACK),
	.NUMBER_STOP_BITS(NUMBER_STOP_BITS),
	.TX_MASSIV_DEEP(TX_MASSIV_DEEP),
	.RX_MASSIV_DEEP(RX_MASSIV_DEEP)
)
TX_RX_MASSIV1
(
	.IN_CLOCK(IN_CLOCK_1),
	.IN_TX_DATA_MASSIV(IN_TX_DATA_MASSIV_1),
	.IN_TX_NUMBER_OF_PACKS_TO_SEND(IN_TX_NUMBER_OF_PACKS_TO_SEND_1),
	.IN_TX_LAUNCH(IN_TX_LAUNCH_1),
	.OUT_TX_ACTIVE(OUT_TX_ACTIVE_1),
	.OUT_TX_DONE(OUT_TX_DONE_1),
	.IN_RX_CLEAR_BUFFER(IN_RX_CLEAR_BUFFER_1),
	.OUT_RX_DATA_MASSIV(OUT_RX_DATA_MASSIV_1),
	.OUT_RX_ERROR(OUT_RX_ERROR_1),
	.OUT_RX_NUM_OF_DATA_PACKS_READY(OUT_RX_NUM_OF_DATA_PACKS_READY_1),
	.TX_PORT(TRANSMIT_1_TO_2),
	.RX_PORT(TRANSMIT_2_TO_1)
);


UART_TX_RX_MASSIV_MODULE
#(
	.UART_BAUD_RATE(UART_BAUD_RATE),
	.CLOCK_FREQUENCY(CLOCK_FREQUENCY),
	.PARITY(PARITY),
	.NUM_OF_DATA_BITS_IN_PACK(NUM_OF_DATA_BITS_IN_PACK),
	.NUMBER_STOP_BITS(NUMBER_STOP_BITS),
	.TX_MASSIV_DEEP(TX_MASSIV_DEEP),
	.RX_MASSIV_DEEP(RX_MASSIV_DEEP)
)
TX_RX_MASSIV2
(
	.IN_CLOCK(IN_CLOCK_2),
	.IN_TX_DATA_MASSIV(IN_TX_DATA_MASSIV_2),
	.IN_TX_NUMBER_OF_PACKS_TO_SEND(IN_TX_NUMBER_OF_PACKS_TO_SEND_1),
	.OUT_TX_ACTIVE(OUT_TX_ACTIVE_2),
	.IN_TX_LAUNCH(IN_TX_LAUNCH_2),
	.OUT_TX_DONE(OUT_TX_DONE_2),
	.IN_RX_CLEAR_BUFFER(IN_RX_CLEAR_BUFFER_2),
	.OUT_RX_DATA_MASSIV(OUT_RX_DATA_MASSIV_2),
	.OUT_RX_ERROR(OUT_RX_ERROR_2),
	.OUT_RX_NUM_OF_DATA_PACKS_READY(OUT_RX_NUM_OF_DATA_PACKS_READY_2),
	.TX_PORT(TRANSMIT_2_TO_1),
	.RX_PORT(TRANSMIT_1_TO_2)
);


always 
	begin
		#(PERIOD_IN_CLOCK_NS/2)
		IN_CLOCK_1=!IN_CLOCK_1;
		IN_CLOCK_2=!IN_CLOCK_2;
	end

	
initial begin
		IN_TX_LAUNCH_1=0;IN_TX_LAUNCH_1=0;
		IN_CLOCK_1=1'b1;IN_CLOCK_2=1'b0;
		IN_TX_DATA_MASSIV_1=0;IN_TX_DATA_MASSIV_2=0;
		#(PERIOD_IN_CLOCK_NS*10)
		IN_TX_DATA_MASSIV_1=16'b0010110000111011;
		IN_TX_DATA_MASSIV_2=16'bZ;
		#(PERIOD_IN_CLOCK_NS*10)
		IN_TX_NUMBER_OF_PACKS_TO_SEND_1=TX_MASSIV_DEEP;
		IN_TX_NUMBER_OF_PACKS_TO_SEND_2=0;
		#(PERIOD_IN_CLOCK_NS*10)
		IN_TX_LAUNCH_1=1;IN_TX_LAUNCH_2=0;
		#(PERIOD_IN_CLOCK_NS*10)
		IN_TX_LAUNCH_1=0;
		
		@(posedge (OUT_RX_NUM_OF_DATA_PACKS_READY_2==2))
		begin
			#(PERIOD_IN_CLOCK_NS*5)
			IN_TX_DATA_MASSIV_2<=OUT_RX_DATA_MASSIV_2[NUM_OF_DATA_BITS_IN_PACK-1:0]+OUT_RX_DATA_MASSIV_2[NUM_OF_DATA_BITS_IN_PACK*2-1:NUM_OF_DATA_BITS_IN_PACK];
			#(PERIOD_IN_CLOCK_NS*10)
			IN_RX_CLEAR_BUFFER_2=1;
			#(PERIOD_IN_CLOCK_NS*10)
			IN_RX_CLEAR_BUFFER_2=0;
			IN_TX_LAUNCH_2=1;
			#(PERIOD_IN_CLOCK_NS*10)
			IN_TX_LAUNCH_2=0;
		end
		@(posedge (OUT_RX_NUM_OF_DATA_PACKS_READY_1==1))
		begin
			#(PERIOD_IN_CLOCK_NS*5)
			IN_TX_DATA_MASSIV_1<=OUT_RX_DATA_MASSIV_1[NUM_OF_DATA_BITS_IN_PACK-1:0]/2;
			#(PERIOD_IN_CLOCK_NS*10)
			IN_RX_CLEAR_BUFFER_1=1;
			#(PERIOD_IN_CLOCK_NS*10)
			IN_RX_CLEAR_BUFFER_1=0;
			IN_TX_LAUNCH_1=1;
			#(PERIOD_IN_CLOCK_NS*10)
			IN_TX_LAUNCH_1=0;
		end
		
	
end
//блок ожидания приемника

endmodule
